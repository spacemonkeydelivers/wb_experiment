`define WB_ADDR_WIDTH 32
`define WB_DATA_WIDTH 16
`define EXT_DATA_WIDTH 16
`define EXT_ADDR_WIDTH 32
`define ITH_BYTE(i) 8*(i+1)-1:8*i
